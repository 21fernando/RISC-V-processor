module csr(
    input clock
);

endmodule