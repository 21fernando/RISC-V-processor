module csr(
    input clock,
    input 
);

endmodule